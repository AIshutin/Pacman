00000000000
00.0...0.00
00..0.0..00
00.0...0.00
0.........0
00000.00000
0..<..a..<0
00.00.00.00
00....c..00
00.00000.00
00000000000

