00000000000000000000
0.0.000000000000<0.0
0.0........<.....0.0
0.0.0.00000000.0.0.0
0...0.00000000.0...0
00.0.....00.....0.00
0...0.00.00.00.0...0
00.0.0........0.0.00
00...0.0.00.0.0...00
00.0.0..<.....0.0.00
00.0.0........0.0.00
00.....0.00.0.....00
00.0.0.....<..0.0.00
00.00.00.00.00.00.00
00.00..0....0..00.00
00.00.00.00.00.00.00
00.00.00.00.00.00.00
00....00.00.00....00
00000.00.00.00.00000
00000000000000000000

