00000
0.0.0
0.<<0
0.0.0
00000

