00000000000
00.00000.00
0<........0
00.00.00<00
00000.00000
0.........0
00.00.00<00
00.00.00.00
0..0<..0..0
00000.00000
00000000000

